module I2S (
	input CLK,
	input RESET,
	input [31:0] Din,
	input LRCLK,
	input SCLK,
	output [31:0] Dout
);

endmodule
